library IEEE;
use IEEE.STD_LOGIC_1164.all;

package DecoderPackage is
Component Decoder is
Port (
        input : in  STD_LOGIC_VECTOR (4 downto 0);
        out0 : out  STD_LOGIC;
        out1 : out  STD_LOGIC;
        out2 : out  STD_LOGIC;
        out3 : out  STD_LOGIC;
        out4 : out  STD_LOGIC;
        out5 : out  STD_LOGIC;
        out6 : out  STD_LOGIC;
        out7 : out  STD_LOGIC;
        out8 : out  STD_LOGIC;
        out9 : out  STD_LOGIC;
        out10 : out  STD_LOGIC;
        out11 : out  STD_LOGIC;
        out12 : out  STD_LOGIC;
        out13 : out  STD_LOGIC;
        out14 : out  STD_LOGIC;
        out15 : out  STD_LOGIC;
        out16 : out  STD_LOGIC;
        out17 : out  STD_LOGIC;
        out18 : out  STD_LOGIC;
        out19 : out  STD_LOGIC;
        out20 : out  STD_LOGIC;
        out21 : out  STD_LOGIC;
        out22 : out  STD_LOGIC;
        out23 : out  STD_LOGIC;
        out24 : out  STD_LOGIC;
        out25 : out  STD_LOGIC;
        out26 : out  STD_LOGIC;
        out27 : out  STD_LOGIC;
        out28 : out  STD_LOGIC;
        out29 : out  STD_LOGIC;
        out30 : out  STD_LOGIC;
        out31 : out  STD_LOGIC
		  );
		  end component;
end DecoderPackage;